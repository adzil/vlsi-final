module processor(iarray, tarray, markin, clk, rst, ena, tout, markout, );



endmodule
